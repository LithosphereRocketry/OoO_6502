// Flag register
`define FLAG_CARRY 0
`define FLAG_ZERO 1
`define FLAG_OVERFLOW 6
`define FLAG_NEGATIVE 7

// Microcode parameters (adjust as microcode gets bigger)
`define UCR_ADDR_WIDTH 9