`timescale 1ns/1ps

module core(
        
    );

endmodule