module middle_end(

);

// arithmetic_pipeline _arith_pipe(

// );

// memory_pipeline _mem_pipe(

// );

// terminate_pipeline _term_pipe(

// );

endmodule