`define FLAG_CARRY 0
`define FLAG_OVERFLOW 6